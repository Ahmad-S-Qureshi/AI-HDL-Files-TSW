module clock_divider (
    input wire clk_in,       // 100 MHz clock input
    input wire reset,        // Synchronous reset
    output reg clk_out       // Divided clock output
);

// Generate the remaining module code using an AI language model, maintaining the specified inputs and outputs.

endmodule
